// You need to generate this component correctly



module imem(address, clock, q);
	input [31:0] address;
	input clock;
	output [31:0] q;
	
//
//	reg [31:0] memory [65535:0];
//
//
//	always @(posedge clock) begin
//		 q <= memory[address];
//	end



endmodule
